library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

package speed_rom is
	constant clk_leds_cnt_len: integer := 22;
	constant adr_len: integer := 5;
	constant num_speeds: integer := 32;
	type rom_speed is array (0 to num_speeds - 1) of unsigned(clk_leds_cnt_len - 1 downto 0);
	constant speeds: rom_speed := (
		0 => "1010100110001010110001",
		1 => "1000001101100101001001",
		2 => "0110101101000010111001",
		3 => "0101101010011110000010",
		4 => "0100111001110001111000",
		5 => "0100010100100111110000",
		6 => "0011110111010101001111",
		7 => "0011011111101001101011",
		8 => "0011001100000110111110",
		9 => "0010111011101101010001",
		10 => "0010101101101111101110",
		11 => "0010100001101101111001",
		12 => "0010010111001111110000",
		13 => "0010001110000011000111",
		14 => "0010000101111001111110",
		15 => "0001111110101001010101",
		16 => "0001111000001000011111",
		17 => "0001110010010000011011",
		18 => "0001101100111011011011",
		19 => "0001101000000100110100",
		20 => "0001100011101000101101",
		21 => "0001011111100011110110",
		22 => "0001011011110011011111",
		23 => "0001011000010101010011",
		24 => "0001010101000111010011",
		25 => "0001010010000111110011",
		26 => "0001001111010101010011",
		27 => "0001001100101110100010",
		28 => "0001001010010010010111",
		29 => "0001000111111111110101",
		30 => "0001000101110110000011",
		31 => "0001000011110100010001");
end package;
