library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

package speed_rom is
	constant clk_leds_cnt_len: integer := 25;
	constant adr_len: integer := 5;
	constant num_speeds: integer := 32;
	type rom_speed is array (0 to num_speeds - 1) of unsigned(clk_leds_cnt_len - 1 downto 0);
	constant speeds: rom_speed := (
		0 => "1101001111101101011110001",
		1 => "1011101011001101010111111",
		2 => "1010010010100111110101111",
		3 => "1001000100100010011110001",
		4 => "0111111111101101100100011",
		5 => "0111000011000010111001011",
		6 => "0110001101100100100010101",
		7 => "0101011110011011111011011",
		8 => "0100110100111000111100111",
		9 => "0100010000010001001101110",
		10 => "0011101111111111010110000",
		11 => "0011010011100010011001010",
		12 => "0010111010011101010101010",
		13 => "0010100100010110100011110",
		14 => "0010010000110111100001000",
		15 => "0001111111101100010100011",
		16 => "0001110000100011011100000",
		17 => "0001100011001101011011000",
		18 => "0001010111011100101010001",
		19 => "0001001101000101001000111",
		20 => "0001000011111100010010001",
		21 => "0000111011111000110001000",
		22 => "0000110100110010010111100",
		23 => "0000101110100001110101110",
		24 => "0000101001000000110011000",
		25 => "0000100100001001100111001",
		26 => "0000011111110111010100010",
		27 => "0000011100000101100010110",
		28 => "0000011000110000011011101",
		29 => "0000010101110100100101101",
		30 => "0000010011001111000000111",
		31 => "0000010000111101000100011");
end package;
