library verilog;
use verilog.vl_types.all;
entity band_pass_direct_vhdl_vlg_vec_tst is
end band_pass_direct_vhdl_vlg_vec_tst;
