library ieee;
use ieee.std_logic_1164.all;

package velocities_rom is
	constant clk_div0_len: integer := 24;
	constant adr_len: integer := 7;
	constant num_velocities: integer := 128;
	type rom_vel is array (0 to num_velocities - 1) of std_logic_vector (clk_div0_len - 1 downto 0);
	constant velocities: rom_vel := (
		0 => "101111101011110000100000",
		1 => "101110110100111011010001",
		2 => "101101111111000101000110",
		3 => "101101001010001100110110",
		4 => "101100010110010001011001",
		5 => "101011100011010001101010",
		6 => "101010110001001100100100",
		7 => "101010000000000001000100",
		8 => "101001001111101110000111",
		9 => "101000100000010010101100",
		10 => "100111110001101101110011",
		11 => "100111000011111110011110",
		12 => "100110010111000011110000",
		13 => "100101101010111100101011",
		14 => "100100111111101000010100",
		15 => "100100010101000101110001",
		16 => "100011101011010100001001",
		17 => "100011000010010010100100",
		18 => "100010011010000000001001",
		19 => "100001110010011100000100",
		20 => "100001001011100101011110",
		21 => "100000100101011011100011",
		22 => "011111111111111101100000",
		23 => "011111011011001010100011",
		24 => "011110110111000001111010",
		25 => "011110010011100010110100",
		26 => "011101110000101100100010",
		27 => "011101001110011110010100",
		28 => "011100101100110111011101",
		29 => "011100001011110111001111",
		30 => "011011101011011100111110",
		31 => "011011001011100111111110",
		32 => "011010101100010111100101",
		33 => "011010001101101011001000",
		34 => "011001101111100001111101",
		35 => "011001010001111011011110",
		36 => "011000110100110111000000",
		37 => "011000011000010011111110",
		38 => "010111111100010001110001",
		39 => "010111100000101111110011",
		40 => "010111000101101101011111",
		41 => "010110101011001010010001",
		42 => "010110010001000101100100",
		43 => "010101110111011110110111",
		44 => "010101011110010101100110",
		45 => "010101000101101001001111",
		46 => "010100101101011001010010",
		47 => "010100010101100101001101",
		48 => "010011111110001100100001",
		49 => "010011100111001110101101",
		50 => "010011010000101011010100",
		51 => "010010111010100001110111",
		52 => "010010100100110001111000",
		53 => "010010001111011010111001",
		54 => "010001111010011100011110",
		55 => "010001100101110110001011",
		56 => "010001010001100111100100",
		57 => "010000111101110000001101",
		58 => "010000101010001111101100",
		59 => "010000010111000101100111",
		60 => "010000000100010001100100",
		61 => "001111110001110011001010",
		62 => "001111011111101001111111",
		63 => "001111001101110101101011",
		64 => "001110111100010101110111",
		65 => "001110101011001010001010",
		66 => "001110011010010010001110",
		67 => "001110001001101101101011",
		68 => "001101111001011100001101",
		69 => "001101101001011101011011",
		70 => "001101011001110001000010",
		71 => "001101001010010110101100",
		72 => "001100111011001110000100",
		73 => "001100101100010110110110",
		74 => "001100011101110000101101",
		75 => "001100001111011011010111",
		76 => "001100000001010110100000",
		77 => "001011110011100001110100",
		78 => "001011100101111101000010",
		79 => "001011011000100111110111",
		80 => "001011001011100010000001",
		81 => "001010111110101011001110",
		82 => "001010110010000011001110",
		83 => "001010100101101001101110",
		84 => "001010011001011110011111",
		85 => "001010001101100001010000",
		86 => "001010000001110001110001",
		87 => "001001110110001111110011",
		88 => "001001101010111011000100",
		89 => "001001011111110011011000",
		90 => "001001010100111000011101",
		91 => "001001001010001010000110",
		92 => "001000111111101000000101",
		93 => "001000110101010010001010",
		94 => "001000101011001000001001",
		95 => "001000100001001001110011",
		96 => "001000010111010110111011",
		97 => "001000001101101111010100",
		98 => "001000000100010010110001",
		99 => "000111111011000001000101",
		100 => "000111110001111010000100",
		101 => "000111101000111101100001",
		102 => "000111100000001011010000",
		103 => "000111010111100011000110",
		104 => "000111001111000100110111",
		105 => "000111000110110000011000",
		106 => "000110111110100101011101",
		107 => "000110110110100011111011",
		108 => "000110101110101011101000",
		109 => "000110100110111100011000",
		110 => "000110011111010110000010",
		111 => "000110010111111000011011",
		112 => "000110010000100011011010",
		113 => "000110001001010110110100",
		114 => "000110000010010010011111",
		115 => "000101111011010110010011",
		116 => "000101110100100010000101",
		117 => "000101101101110101101101",
		118 => "000101100111010001000001",
		119 => "000101100000110011111010",
		120 => "000101011010011110001101",
		121 => "000101010100001111110011",
		122 => "000101001110001000100011",
		123 => "000101001000001000010101",
		124 => "000101000010001111000000",
		125 => "000100111100011100011110",
		126 => "000100110110110000100101",
		127 => "000100110001001011010000");
end package;
