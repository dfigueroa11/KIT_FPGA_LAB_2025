library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

package speed_rom is
	constant clk_leds_cnt_len: integer := 25;
	constant adr_len: integer := 5;
	constant num_speeds: integer := 32;
	type rom_speed is array (0 to num_speeds - 1) of unsigned(clk_leds_cnt_len - 1 downto 0);
	constant speeds: rom_speed := (
		0 => "1101001111101101011110001",
		1 => "0101001000011111001110000",
		2 => "0011001011101101101001111",
		3 => "0010010011101000101000110",
		4 => "0001110011110001000100001",
		5 => "0001011111001101101011111",
		6 => "0001010000110110111100100",
		7 => "0001000110010000111100100",
		8 => "0000111110001000000001011",
		9 => "0000110111101011010000011",
		10 => "0000110010011100001000100",
		11 => "0000101110000110101000001",
		12 => "0000101010011101000011100",
		13 => "0000100111010101110000000",
		14 => "0000100100101001101011111",
		15 => "0000100010010011101000101",
		16 => "0000100000001111101000010",
		17 => "0000011110011010100110000",
		18 => "0000011100110010000111110",
		19 => "0000011011010100010010101",
		20 => "0000011001111111100011101",
		21 => "0000011000110010101010000",
		22 => "0000010111101100100011011",
		23 => "0000010110101100011000011",
		24 => "0000010101110001011010110",
		25 => "0000010100111011000011110",
		26 => "0000010100001000110001111",
		27 => "0000010011011010001000111",
		28 => "0000010010101110110000100",
		29 => "0000010010000110010011011",
		30 => "0000010001100000011111011",
		31 => "0000010000111101000100011");
end package;
