library verilog;
use verilog.vl_types.all;
entity high_pass_transposed_graph_vlg_vec_tst is
end high_pass_transposed_graph_vlg_vec_tst;
