LIBRARY IEEE;
USE IEEE.std_logic_1164.ALL;

PACKAGE my_pkg IS
    SUBTYPE bit4 IS std_logic_vector(7 downto 0);
END my_pkg;
