library verilog;
use verilog.vl_types.all;
entity band_stop_transposed_vhdl_vlg_vec_tst is
end band_stop_transposed_vhdl_vlg_vec_tst;
