library verilog;
use verilog.vl_types.all;
entity low_pass_direct_graph_vlg_vec_tst is
end low_pass_direct_graph_vlg_vec_tst;
