library ieee;
use ieee.std_logic_1164.all;

package speed_rom is
	constant clk_div0_len: integer := 23;
	constant adr_len: integer := 8;
	constant num_speeds: integer := 256;
	type rom_speed is array (0 to num_speeds - 1) of std_logic_vector (clk_div0_len - 1 downto 0);
	constant speeds: rom_speed := (
		0 => "10111110101111000010000",
		1 => "10111000001110111000011",
		2 => "10110010001010001011000",
		3 => "10101100011110010001011",
		4 => "10100111001000111000100",
		5 => "10100010000111111110011",
		6 => "10011101011001110000110",
		7 => "10011000111100101010000",
		8 => "10010100101111001111101",
		9 => "10010000110000010000111",
		10 => "10001100111110100101101",
		11 => "10001001011001001100110",
		12 => "10000101111111001011111",
		13 => "10000010101111101110010",
		14 => "01111111101010000011110",
		15 => "01111100101101100001010",
		16 => "01111001111001011111000",
		17 => "01110111001101011001001",
		18 => "01110100101000101110110",
		19 => "01110010001011000001101",
		20 => "01101111110011110110001",
		21 => "01101101100010110010111",
		22 => "01101011010111100000011",
		23 => "01101001010001101001011",
		24 => "01100111010000111001101",
		25 => "01100101010100111111000",
		26 => "01100011011101101000010",
		27 => "01100001101010100101101",
		28 => "01011111111011101000011",
		29 => "01011110010000100010110",
		30 => "01011100101001001000010",
		31 => "01011011000101001100110",
		32 => "01011001100100100101010",
		33 => "01011000000111000111100",
		34 => "01010110101100101001101",
		35 => "01010101010101000010100",
		36 => "01010100000000001001110",
		37 => "01010010101101110111011",
		38 => "01010001011110000011101",
		39 => "01010000010000100111110",
		40 => "01001111000101011100111",
		41 => "01001101111100011100110",
		42 => "01001100110101100001100",
		43 => "01001011110000100101100",
		44 => "01001010101101100011100",
		45 => "01001001101100010110100",
		46 => "01001000101100111001110",
		47 => "01000111101111001000111",
		48 => "01000110110010111111100",
		49 => "01000101111000011001110",
		50 => "01000100111111010011110",
		51 => "01000100000111101001110",
		52 => "01000011010001011000100",
		53 => "01000010011100011100110",
		54 => "01000001101000110011001",
		55 => "01000000110110011000111",
		56 => "01000000000101001011010",
		57 => "00111111010101000111011",
		58 => "00111110100110001010110",
		59 => "00111101111000010010111",
		60 => "00111101001011011101100",
		61 => "00111100011111101000100",
		62 => "00111011110100110001100",
		63 => "00111011001010110110100",
		64 => "00111010100001110101110",
		65 => "00111001111001101101001",
		66 => "00111001010010011011000",
		67 => "00111000101011111101101",
		68 => "00111000000110010011011",
		69 => "00110111100001011010101",
		70 => "00110110111101010001111",
		71 => "00110110011001110111110",
		72 => "00110101110111001010110",
		73 => "00110101010101001001100",
		74 => "00110100110011110011000",
		75 => "00110100010011000101101",
		76 => "00110011110011000000100",
		77 => "00110011010011100010010",
		78 => "00110010110100101010000",
		79 => "00110010010110010110100",
		80 => "00110001111000100110111",
		81 => "00110001011011011010000",
		82 => "00110000111110101111000",
		83 => "00110000100010100101000",
		84 => "00110000000110111011001",
		85 => "00101111101011110000100",
		86 => "00101111010001000100001",
		87 => "00101110110110110101100",
		88 => "00101110011101000011110",
		89 => "00101110000011101110000",
		90 => "00101101101010110011110",
		91 => "00101101010010010100010",
		92 => "00101100111010001110110",
		93 => "00101100100010100010110",
		94 => "00101100001011001111011",
		95 => "00101011110100010100010",
		96 => "00101011011101110000110",
		97 => "00101011000111100100010",
		98 => "00101010110001101110011",
		99 => "00101010011100001110010",
		100 => "00101010000111000011110",
		101 => "00101001110010001110001",
		102 => "00101001011101101100111",
		103 => "00101001001001011111110",
		104 => "00101000110101100110001",
		105 => "00101000100001111111100",
		106 => "00101000001110101011110",
		107 => "00100111111011101010001",
		108 => "00100111101000111010011",
		109 => "00100111010110011100001",
		110 => "00100111000100001111000",
		111 => "00100110110010010010101",
		112 => "00100110100000100110100",
		113 => "00100110001111001010100",
		114 => "00100101111101111110001",
		115 => "00100101101101000001001",
		116 => "00100101011100010011001",
		117 => "00100101001011110011111",
		118 => "00100100111011100011000",
		119 => "00100100101011100000011",
		120 => "00100100011011101011100",
		121 => "00100100001100000100001",
		122 => "00100011111100101010001",
		123 => "00100011101101011101010",
		124 => "00100011011110011101000",
		125 => "00100011001111101001011",
		126 => "00100011000001000010000",
		127 => "00100010110010100110101",
		128 => "00100010100100010111001",
		129 => "00100010010110010011001",
		130 => "00100010001000011010101",
		131 => "00100001111010101101001",
		132 => "00100001101101001010101",
		133 => "00100001011111110010111",
		134 => "00100001010010100101110",
		135 => "00100001000101100010111",
		136 => "00100000111000101010010",
		137 => "00100000101011111011100",
		138 => "00100000011111010110101",
		139 => "00100000010010111011010",
		140 => "00100000000110101001100",
		141 => "00011111111010100000111",
		142 => "00011111101110100001100",
		143 => "00011111100010101011000",
		144 => "00011111010110111101010",
		145 => "00011111001011011000010",
		146 => "00011110111111111011110",
		147 => "00011110110100100111100",
		148 => "00011110101001011011101",
		149 => "00011110011110010111110",
		150 => "00011110010011011011110",
		151 => "00011110001000100111101",
		152 => "00011101111101111011001",
		153 => "00011101110011010110010",
		154 => "00011101101000111000110",
		155 => "00011101011110100010101",
		156 => "00011101010100010011101",
		157 => "00011101001010001011101",
		158 => "00011101000000001010101",
		159 => "00011100110110010000100",
		160 => "00011100101100011101001",
		161 => "00011100100010110000011",
		162 => "00011100011001001010001",
		163 => "00011100001111101010010",
		164 => "00011100000110010000110",
		165 => "00011011111100111101100",
		166 => "00011011110011110000010",
		167 => "00011011101010101001001",
		168 => "00011011100001101000000",
		169 => "00011011011000101100101",
		170 => "00011011001111110111001",
		171 => "00011011000111000111001",
		172 => "00011010111110011100111",
		173 => "00011010110101111000000",
		174 => "00011010101101011000101",
		175 => "00011010100100111110101",
		176 => "00011010011100101001111",
		177 => "00011010010100011010010",
		178 => "00011010001100001111111",
		179 => "00011010000100001010011",
		180 => "00011001111100001010000",
		181 => "00011001110100001110011",
		182 => "00011001101100010111101",
		183 => "00011001100100100101101",
		184 => "00011001011100111000011",
		185 => "00011001010101001111110",
		186 => "00011001001101101011101",
		187 => "00011001000110001100000",
		188 => "00011000111110110000111",
		189 => "00011000110111011010000",
		190 => "00011000110000000111100",
		191 => "00011000101000111001010",
		192 => "00011000100001101111010",
		193 => "00011000011010101001011",
		194 => "00011000010011100111100",
		195 => "00011000001100101001110",
		196 => "00011000000101101111111",
		197 => "00010111111110111010000",
		198 => "00010111111000001000000",
		199 => "00010111110001011001110",
		200 => "00010111101010101111011",
		201 => "00010111100100001000101",
		202 => "00010111011101100101101",
		203 => "00010111010111000110001",
		204 => "00010111010000101010011",
		205 => "00010111001010010010000",
		206 => "00010111000011111101001",
		207 => "00010110111101101011110",
		208 => "00010110110111011101110",
		209 => "00010110110001010011001",
		210 => "00010110101011001011110",
		211 => "00010110100101000111110",
		212 => "00010110011111000110111",
		213 => "00010110011001001001010",
		214 => "00010110010011001110110",
		215 => "00010110001101010111011",
		216 => "00010110000111100011001",
		217 => "00010110000001110001111",
		218 => "00010101111100000011100",
		219 => "00010101110110011000010",
		220 => "00010101110000101111111",
		221 => "00010101101011001010011",
		222 => "00010101100101100111110",
		223 => "00010101100000000111111",
		224 => "00010101011010101010111",
		225 => "00010101010101010000101",
		226 => "00010101001111111001000",
		227 => "00010101001010100100001",
		228 => "00010101000101010010000",
		229 => "00010101000000000010011",
		230 => "00010100111010110101011",
		231 => "00010100110101101011000",
		232 => "00010100110000100011001",
		233 => "00010100101011011101110",
		234 => "00010100100110011010111",
		235 => "00010100100001011010100",
		236 => "00010100011100011100100",
		237 => "00010100010111100000111",
		238 => "00010100010010100111101",
		239 => "00010100001101110000110",
		240 => "00010100001000111100001",
		241 => "00010100000100001001111",
		242 => "00010011111111011001111",
		243 => "00010011111010101100001",
		244 => "00010011110110000000100",
		245 => "00010011110001010111001",
		246 => "00010011101100110000000",
		247 => "00010011101000001010111",
		248 => "00010011100011101000000",
		249 => "00010011011111000111001",
		250 => "00010011011010101000011",
		251 => "00010011010110001011101",
		252 => "00010011010001110001000",
		253 => "00010011001101011000011",
		254 => "00010011001001000001101",
		255 => "00010011000100101101000");
end package;
